`timescale 1ns / 1ps

module OR(
input x,y,
output o
);

assign o = x|y;


endmodule
