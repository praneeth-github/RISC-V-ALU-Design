`timescale 1ns / 1ps
module OR(
	input A,B,
	output O
	);
	
	assign O = A | B;

endmodule
