`timescale 1ns / 1ps

module AND(
input x,y,
output o
);

assign o = x & y;

endmodule
