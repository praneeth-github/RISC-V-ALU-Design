`timescale 1ns / 1ps
module AND(
	input A,B,
	output O
	);
	
	assign O = A & B;

endmodule